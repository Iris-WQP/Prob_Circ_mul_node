`define DW 16     //BF16
`define Tin 8
`define Tout 4
`define bram_depth_in 2048
`define log2_bram_depth_in 11
`define bram_width_in `DW*`Tin //128