`define DW 16     //BF16